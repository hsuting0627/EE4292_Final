module top(
    input clk,
    input rst_n,
    input enable,
    input [512-1:0] data_read,
    output [11-1:0] sram_raddr,
    output [11-1:0] sram_waddr,
    output [512-1:0] data_write,
    output  [10:0]  q11, q12, q13, q14, q15, q16, q17, q18, q21, q22, q23, q24,
    output  [10:0]  q25, q26, q27, q28, q31, q32, q33, q34, q35, q36, q37, q38,
    output  [10:0]  q41, q42, q43, q44, q45, q46, q47, q48, q51, q52, q53, q54,
    output  [10:0]  q55, q56, q57, q58, q61, q62, q63, q64, q65, q66, q67, q68,
    output  [10:0]  q71, q72, q73, q74, q75, q76, q77, q78, q81, q82, q83, q84,
    output  [10:0]  q85, q86, q87, q88,
    output wen,
    output valid
);
//====== Control Unit =======
wire enable_rgb2ycbcr;
wire valid_rgb2ycbcr;
wire enable_dct;
wire enable_quan;
wire valid_dct;
wire valid_quan;
wire [10:0] sram_raddr_dct, sram_raddr_rgb2ycbcr;
assign sram_raddr = enable_rgb2ycbcr ? sram_raddr_rgb2ycbcr : sram_raddr_dct;
// === variable here is for testing dat format and can be deleted if you have other purposes.
    wire signed [11-1:0] dct00, dct01, dct02, dct03, dct04, dct05, dct06, dct07;
    wire signed [11-1:0] dct10, dct11, dct12, dct13, dct14, dct15, dct16, dct17;
    wire signed [11-1:0] dct20, dct21, dct22, dct23, dct24, dct25, dct26, dct27;
    wire signed [11-1:0] dct30, dct31, dct32, dct33, dct34, dct35, dct36, dct37;
    wire signed [11-1:0] dct40, dct41, dct42, dct43, dct44, dct45, dct46, dct47;
    wire signed [11-1:0] dct50, dct51, dct52, dct53, dct54, dct55, dct56, dct57;
    wire signed [11-1:0] dct60, dct61, dct62, dct63, dct64, dct65, dct66, dct67;
    wire signed [11-1:0] dct70, dct71, dct72, dct73, dct74, dct75, dct76, dct77;
//===========================================================================================

// controller here is for rgb2ycbcr and dct.
// the valid_dct means that the data can be quantized !
// the done_dct is for testing here for rgb2ycbcr, and can be removed if you want to add quantization module.
// add control signal here to control the quantization and huffman table !
// good luck! (I need to study RFIC q_q)

// wire  [10:0]  q11, q12, q13, q14, q15, q16, q17, q18, q21, q22, q23, q24;
// wire  [10:0]  q25, q26, q27, q28, q31, q32, q33, q34, q35, q36, q37, q38;
// wire  [10:0]  q41, q42, q43, q44, q45, q46, q47, q48, q51, q52, q53, q54;
// wire  [10:0]  q55, q56, q57, q58, q61, q62, q63, q64, q65, q66, q67, q68;
// wire  [10:0]  q71, q72, q73, q74, q75, q76, q77, q78, q81, q82, q83, q84;
// wire  [10:0]  q85, q86, q87, q88;

controller controller (
    .clk(clk),
    .rst_n(rst_n),
    .enable(enable),
    .enable_rgb2ycbcr(enable_rgb2ycbcr),
    .valid_rgb2ycbcr(valid_rgb2ycbcr),
    .enable_dct(enable_dct),
    .enable_quan(enable_quan),
    .valid_dct(valid_dct),
    .valid_quan(valid_quan),
    .valid(valid)//
);

rgb2ycbcr_2d rgb2ycbcr_2d (
    .clk(clk),
    .rst_n(rst_n),
    .enable(enable_rgb2ycbcr),
    .data_read(data_read), 
    .sram_raddr(sram_raddr_rgb2ycbcr),
    .sram_waddr(sram_waddr),
    .data_write(data_write), 
    .wen(wen),
    .valid(valid_rgb2ycbcr)
);

dct_2d dct_2d (
    .clk(clk),
    .rst_n(rst_n),
    .enable(enable_dct),
    .data_read(data_read),
    .sram_raddr(sram_raddr_dct),
    .valid(valid_dct),
    // .done(done_dct),
    .dct00(dct00),
    .dct01(dct01),
    .dct02(dct02),
    .dct03(dct03),
    .dct04(dct04),
    .dct05(dct05),
    .dct06(dct06),
    .dct07(dct07),
    .dct10(dct10),
    .dct11(dct11),
    .dct12(dct12),
    .dct13(dct13),
    .dct14(dct14),
    .dct15(dct15),
    .dct16(dct16),
    .dct17(dct17),
    .dct20(dct20),
    .dct21(dct21),
    .dct22(dct22),
    .dct23(dct23),
    .dct24(dct24),
    .dct25(dct25),
    .dct26(dct26),
    .dct27(dct27),
    .dct30(dct30),
    .dct31(dct31),
    .dct32(dct32),
    .dct33(dct33),
    .dct34(dct34),
    .dct35(dct35),
    .dct36(dct36),
    .dct37(dct37),
    .dct40(dct40),
    .dct41(dct41),
    .dct42(dct42),
    .dct43(dct43),
    .dct44(dct44),
    .dct45(dct45),
    .dct46(dct46),
    .dct47(dct47),
    .dct50(dct50),
    .dct51(dct51),
    .dct52(dct52),
    .dct53(dct53),
    .dct54(dct54),
    .dct55(dct55),
    .dct56(dct56),
    .dct57(dct57),
    .dct60(dct60),
    .dct61(dct61),
    .dct62(dct62),
    .dct63(dct63),
    .dct64(dct64),
    .dct65(dct65),
    .dct66(dct66),
    .dct67(dct67),
    .dct70(dct70),
    .dct71(dct71),
    .dct72(dct72),
    .dct73(dct73),
    .dct74(dct74),
    .dct75(dct75),
    .dct76(dct76),
    .dct77(dct77)
);

// === variable here is for testing dat format and can be deleted if you have other purposes.
// wire [704-1:0] dct;
// assign dct = {dct00, dct01, dct02, dct03, dct04, dct05, dct06, dct07, dct10, dct11, dct12, dct13, dct14, dct15, dct16, dct17, dct20, dct21, dct22, dct23, dct24, dct25, dct26, dct27, dct30, dct31, dct32, dct33, dct34, dct35, dct36, dct37, dct40, dct41, dct42, dct43, dct44, dct45, dct46, dct47, dct50, dct51, dct52, dct53, dct54, dct55, dct56, dct57, dct60, dct61, dct62, dct63, dct64, dct65, dct66, dct67, dct70, dct71, dct72, dct73, dct74, dct75, dct76, dct77};
//===========================================================================================

quantizer q1(
    .clk(clk), 
    .srst_n(rst_n),
    .enable(enable_quan),
    .mode(1'b0),
    .dct11(dct00),
    .dct12(dct01),
    .dct13(dct02),
    .dct14(dct03),
    .dct15(dct04),
    .dct16(dct05),
    .dct17(dct06),
    .dct18(dct07),
    .dct21(dct10),
    .dct22(dct11),
    .dct23(dct12),
    .dct24(dct13),
    .dct25(dct14),
    .dct26(dct15),
    .dct27(dct16),
    .dct28(dct17),
    .dct31(dct20),
    .dct32(dct21),
    .dct33(dct22),
    .dct34(dct23),
    .dct35(dct24),
    .dct36(dct25),
    .dct37(dct26),
    .dct38(dct27),
    .dct41(dct30),
    .dct42(dct31),
    .dct43(dct32),
    .dct44(dct33),
    .dct45(dct34),
    .dct46(dct35),
    .dct47(dct36),
    .dct48(dct37),
    .dct51(dct40),
    .dct52(dct41),
    .dct53(dct42),
    .dct54(dct43),
    .dct55(dct44),
    .dct56(dct45),
    .dct57(dct46),
    .dct58(dct47),
    .dct61(dct50),
    .dct62(dct51),
    .dct63(dct52),
    .dct64(dct53),
    .dct65(dct54),
    .dct66(dct55),
    .dct67(dct56),
    .dct68(dct57),
    .dct71(dct60),
    .dct72(dct61),
    .dct73(dct62),
    .dct74(dct63),
    .dct75(dct64),
    .dct76(dct65),
    .dct77(dct66),
    .dct78(dct67),
    .dct81(dct70),
    .dct82(dct71),
    .dct83(dct72),
    .dct84(dct73),
    .dct85(dct74),
    .dct86(dct75),
    .dct87(dct76),
    .dct88(dct77),
    .q11(q11),
    .q12(q12),
    .q13(q13),
    .q14(q14),
    .q15(q15),
    .q16(q16),
    .q17(q17),
    .q18(q18),
    .q21(q21),
    .q22(q22),
    .q23(q23),
    .q24(q24),
    .q25(q25),
    .q26(q26),
    .q27(q27),
    .q28(q28),
    .q31(q31),
    .q32(q32),
    .q33(q33),
    .q34(q34),
    .q35(q35),
    .q36(q36),
    .q37(q37),
    .q38(q38),
    .q41(q41),
    .q42(q42),
    .q43(q43),
    .q44(q44),
    .q45(q45),
    .q46(q46),
    .q47(q47),
    .q48(q48),
    .q51(q51),
    .q52(q52),
    .q53(q53),
    .q54(q54),
    .q55(q55),
    .q56(q56),
    .q57(q57),
    .q58(q58),
    .q61(q61),
    .q62(q62),
    .q63(q63),
    .q64(q64),
    .q65(q65),
    .q66(q66),
    .q67(q67),
    .q68(q68),
    .q71(q71),
    .q72(q72),
    .q73(q73),
    .q74(q74),
    .q75(q75),
    .q76(q76),
    .q77(q77),
    .q78(q78),
    .q81(q81),
    .q82(q82),
    .q83(q83),
    .q84(q84),
    .q85(q85),
    .q86(q86),
    .q87(q87),
    .q88(q88),
    .vaild(valid_quan)
);

// RLC e1(
// 	.clk(clk), 
//     .srst_n(srst_n),
//     .q11(q11),
//     .q12(q12),
//     .q13(q13),
//     .q14(q14),
//     .q15(q15),
//     .q16(q16),
//     .q17(q17),
//     .q18(q18),
//     .q21(q21),
//     .q22(q22),
//     .q23(q23),
//     .q24(q24),
//     .q25(q25),
//     .q26(q26),
//     .q27(q27),
//     .q28(q28),
//     .q31(q31),
//     .q32(q32),
//     .q33(q33),
//     .q34(q34),
//     .q35(q35),
//     .q36(q36),
//     .q37(q37),
//     .q38(q38),
//     .q41(q41),
//     .q42(q42),
//     .q43(q43),
//     .q44(q44),
//     .q45(q45),
//     .q46(q46),
//     .q47(q47),
//     .q48(q48),
//     .q51(q51),
//     .q52(q52),
//     .q53(q53),
//     .q54(q54),
//     .q55(q55),
//     .q56(q56),
//     .q57(q57),
//     .q58(q58),
//     .q61(q61),
//     .q62(q62),
//     .q63(q63),
//     .q64(q64),
//     .q65(q65),
//     .q66(q66),
//     .q67(q67),
//     .q68(q68),
//     .q71(q71),
//     .q72(q72),
//     .q73(q73),
//     .q74(q74),
//     .q75(q75),
//     .q76(q76),
//     .q77(q77),
//     .q78(q78),
//     .q81(q81),
//     .q82(q82),
//     .q83(q83),
//     .q84(q84),
//     .q85(q85),
//     .q86(q86),
//     .q87(q87),
//     .q88(q88),
//     .enable(vaild_1),
// 	.DC_reg(DC),
// 	.R_reg(R),
// 	.L_reg(L),
// 	.F_reg(F),
// 	.sram_waddr(sram_waddr),
// 	.sram_wdata(sram_wdata),
// 	.wen(wen),
// 	.vaild(vaild)
// );

// always @* begin
//     data_out = {q11, q12, q13, q14, q15, q16, q17, q18, q21, q22, q23, q24, q25, q26, q27, q28, q31, q32, q33, q34, q35, q36, q37, q38, q41, q42, q43, q44, q45, q46, q47, q48, q51, q52, q53, q54, q55, q56, q57, q58, q61, q62, q63, q64, q65, q66, q67, q68, q71, q72, q73, q74, q75, q76, q77, q78, q81, q82, q83, q84, q85, q86, q87, q88};
// end
endmodule