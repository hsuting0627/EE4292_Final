`define N 10
`define M 12

module top(
	input		clk,
	input		rst_n,
	input		enable,
	input		mode,

    output [11-1:0] sramA_raddr,
    input [512-1:0] sramA_rdata,
    output [11-1:0] sramA_waddr,
    output [512-1:0] sramA_wdata,
    output sramA_wen,

	// output  [`N:0] DC,
	// output  [24-1:0] R,
	// output  [32-1:0] L,
	// output  [32-1:0] F,

    output  [11-1:0] sramB_raddr,
    input  [99-1:0] sramB_rdata,
	output  [11-1:0] sramB_waddr,
    output  [99-1:0] sramB_wdata,
    output sramB_wen,

    output [5-1:0] code_length1,
    output [5-1:0] code_length2,
    output [5-1:0] code_length3,
    output [5-1:0] code_length4,
    output [5-1:0] code_length5,
    output [5-1:0] code_length6,
    output [5-1:0] code_length7,
    output [5-1:0] code_length8,
    output [32-1:0] code_out1,
    output [32-1:0] code_out2,
    output [32-1:0] code_out3,
    output [32-1:0] code_out4,
    output [32-1:0] code_out5,
    output [32-1:0] code_out6,
    output [32-1:0] code_out7,
    output [32-1:0] code_out8,
    output [5-1:0] code_length_DC,
    output [20-1:0] code_out_DC,
    output [5-1:0] code_length_table,
    output [32-1:0] code_out_table,
    output out_valid

);
//====== Control Unit =======
wire enable_rgb2ycbcr;
wire enable_dct;
wire enable_quan;
wire enable_RLC;
wire enable_huffman;
wire valid_rgb2ycbcr;
wire valid_dct;
wire valid_quan;
wire valid_RLC;
wire valid_huffman;

wire [10:0] sram_raddr_dct, sram_raddr_rgb2ycbcr;
assign sramA_raddr = valid_rgb2ycbcr ? sram_raddr_dct : sram_raddr_rgb2ycbcr;

wire  [`N:0]  q11, q12, q13, q14, q15, q16, q17, q18, q21, q22, q23, q24;
wire  [`N:0]  q25, q26, q27, q28, q31, q32, q33, q34, q35, q36, q37, q38;
wire  [`N:0]  q41, q42, q43, q44, q45, q46, q47, q48, q51, q52, q53, q54;
wire  [`N:0]  q55, q56, q57, q58, q61, q62, q63, q64, q65, q66, q67, q68;
wire  [`N:0]  q71, q72, q73, q74, q75, q76, q77, q78, q81, q82, q83, q84;
wire  [`N:0]  q85, q86, q87, q88;
    wire signed [11-1:0] dct00, dct01, dct02, dct03, dct04, dct05, dct06, dct07;
    wire signed [11-1:0] dct10, dct11, dct12, dct13, dct14, dct15, dct16, dct17;
    wire signed [11-1:0] dct20, dct21, dct22, dct23, dct24, dct25, dct26, dct27;
    wire signed [11-1:0] dct30, dct31, dct32, dct33, dct34, dct35, dct36, dct37;
    wire signed [11-1:0] dct40, dct41, dct42, dct43, dct44, dct45, dct46, dct47;
    wire signed [11-1:0] dct50, dct51, dct52, dct53, dct54, dct55, dct56, dct57;
    wire signed [11-1:0] dct60, dct61, dct62, dct63, dct64, dct65, dct66, dct67;
    wire signed [11-1:0] dct70, dct71, dct72, dct73, dct74, dct75, dct76, dct77;
rgb2ycbcr_2d rgb2ycbcr_2d (
    .clk(clk),
    .rst_n(rst_n),
    .enable(enable),
    .data_read(sramA_rdata), 
    .sram_raddr(sram_raddr_rgb2ycbcr),
    .sram_waddr(sramA_waddr),
    .data_write(sramA_wdata), 
    .wen(sramA_wen),
    .valid(valid_rgb2ycbcr)
);

dct_2d dct(
    .clk(clk),
    .rst_n(rst_n),
    .enable(valid_rgb2ycbcr), //
    .data_read(sramA_rdata),
    .sram_raddr(sram_raddr_dct),
    .valid(valid_dct),
    // .done(done_dct),
    .dct00(dct00),
    .dct01(dct01),
    .dct02(dct02),
    .dct03(dct03),
    .dct04(dct04),
    .dct05(dct05),
    .dct06(dct06),
    .dct07(dct07),
    .dct10(dct10),
    .dct11(dct11),
    .dct12(dct12),
    .dct13(dct13),
    .dct14(dct14),
    .dct15(dct15),
    .dct16(dct16),
    .dct17(dct17),
    .dct20(dct20),
    .dct21(dct21),
    .dct22(dct22),
    .dct23(dct23),
    .dct24(dct24),
    .dct25(dct25),
    .dct26(dct26),
    .dct27(dct27),
    .dct30(dct30),
    .dct31(dct31),
    .dct32(dct32),
    .dct33(dct33),
    .dct34(dct34),
    .dct35(dct35),
    .dct36(dct36),
    .dct37(dct37),
    .dct40(dct40),
    .dct41(dct41),
    .dct42(dct42),
    .dct43(dct43),
    .dct44(dct44),
    .dct45(dct45),
    .dct46(dct46),
    .dct47(dct47),
    .dct50(dct50),
    .dct51(dct51),
    .dct52(dct52),
    .dct53(dct53),
    .dct54(dct54),
    .dct55(dct55),
    .dct56(dct56),
    .dct57(dct57),
    .dct60(dct60),
    .dct61(dct61),
    .dct62(dct62),
    .dct63(dct63),
    .dct64(dct64),
    .dct65(dct65),
    .dct66(dct66),
    .dct67(dct67),
    .dct70(dct70),
    .dct71(dct71),
    .dct72(dct72),
    .dct73(dct73),
    .dct74(dct74),
    .dct75(dct75),
    .dct76(dct76),
    .dct77(dct77)
);
wire [704-1:0] dct_data;
assign dct_data = {dct00, dct01, dct02, dct03, dct04, dct05, dct06, dct07, dct10, dct11, dct12, dct13, dct14, dct15, dct16, dct17, dct20, dct21, dct22, dct23, dct24, dct25, dct26, dct27, dct30, dct31, dct32, dct33, dct34, dct35, dct36, dct37, dct40, dct41, dct42, dct43, dct44, dct45, dct46, dct47, dct50, dct51, dct52, dct53, dct54, dct55, dct56, dct57, dct60, dct61, dct62, dct63, dct64, dct65, dct66, dct67, dct70, dct71, dct72, dct73, dct74, dct75, dct76, dct77};
quantizer q1(
    .clk(clk), 
    .srst_n(rst_n),
    .enable(valid_dct),
    .mode(mode),
    .dct11(dct00),
    .dct12(dct01),
    .dct13(dct02),
    .dct14(dct03),
    .dct15(dct04),
    .dct16(dct05),
    .dct17(dct06),
    .dct18(dct07),
    .dct21(dct10),
    .dct22(dct11),
    .dct23(dct12),
    .dct24(dct13),
    .dct25(dct14),
    .dct26(dct15),
    .dct27(dct16),
    .dct28(dct17),
    .dct31(dct20),
    .dct32(dct21),
    .dct33(dct22),
    .dct34(dct23),
    .dct35(dct24),
    .dct36(dct25),
    .dct37(dct26),
    .dct38(dct27),
    .dct41(dct30),
    .dct42(dct31),
    .dct43(dct32),
    .dct44(dct33),
    .dct45(dct34),
    .dct46(dct35),
    .dct47(dct36),
    .dct48(dct37),
    .dct51(dct40),
    .dct52(dct41),
    .dct53(dct42),
    .dct54(dct43),
    .dct55(dct44),
    .dct56(dct45),
    .dct57(dct46),
    .dct58(dct47),
    .dct61(dct50),
    .dct62(dct51),
    .dct63(dct52),
    .dct64(dct53),
    .dct65(dct54),
    .dct66(dct55),
    .dct67(dct56),
    .dct68(dct57),
    .dct71(dct60),
    .dct72(dct61),
    .dct73(dct62),
    .dct74(dct63),
    .dct75(dct64),
    .dct76(dct65),
    .dct77(dct66),
    .dct78(dct67),
    .dct81(dct70),
    .dct82(dct71),
    .dct83(dct72),
    .dct84(dct73),
    .dct85(dct74),
    .dct86(dct75),
    .dct87(dct76),
    .dct88(dct77),
    .q11(q11),
    .q12(q12),
    .q13(q13),
    .q14(q14),
    .q15(q15),
    .q16(q16),
    .q17(q17),
    .q18(q18),
    .q21(q21),
    .q22(q22),
    .q23(q23),
    .q24(q24),
    .q25(q25),
    .q26(q26),
    .q27(q27),
    .q28(q28),
    .q31(q31),
    .q32(q32),
    .q33(q33),
    .q34(q34),
    .q35(q35),
    .q36(q36),
    .q37(q37),
    .q38(q38),
    .q41(q41),
    .q42(q42),
    .q43(q43),
    .q44(q44),
    .q45(q45),
    .q46(q46),
    .q47(q47),
    .q48(q48),
    .q51(q51),
    .q52(q52),
    .q53(q53),
    .q54(q54),
    .q55(q55),
    .q56(q56),
    .q57(q57),
    .q58(q58),
    .q61(q61),
    .q62(q62),
    .q63(q63),
    .q64(q64),
    .q65(q65),
    .q66(q66),
    .q67(q67),
    .q68(q68),
    .q71(q71),
    .q72(q72),
    .q73(q73),
    .q74(q74),
    .q75(q75),
    .q76(q76),
    .q77(q77),
    .q78(q78),
    .q81(q81),
    .q82(q82),
    .q83(q83),
    .q84(q84),
    .q85(q85),
    .q86(q86),
    .q87(q87),
    .q88(q88),
    .valid(valid_quan)
);

RLC e1(
	.clk(clk), 
    .srst_n(rst_n),
    .q11(q11),
    .q12(q12),
    .q13(q13),
    .q14(q14),
    .q15(q15),
    .q16(q16),
    .q17(q17),
    .q18(q18),
    .q21(q21),
    .q22(q22),
    .q23(q23),
    .q24(q24),
    .q25(q25),
    .q26(q26),
    .q27(q27),
    .q28(q28),
    .q31(q31),
    .q32(q32),
    .q33(q33),
    .q34(q34),
    .q35(q35),
    .q36(q36),
    .q37(q37),
    .q38(q38),
    .q41(q41),
    .q42(q42),
    .q43(q43),
    .q44(q44),
    .q45(q45),
    .q46(q46),
    .q47(q47),
    .q48(q48),
    .q51(q51),
    .q52(q52),
    .q53(q53),
    .q54(q54),
    .q55(q55),
    .q56(q56),
    .q57(q57),
    .q58(q58),
    .q61(q61),
    .q62(q62),
    .q63(q63),
    .q64(q64),
    .q65(q65),
    .q66(q66),
    .q67(q67),
    .q68(q68),
    .q71(q71),
    .q72(q72),
    .q73(q73),
    .q74(q74),
    .q75(q75),
    .q76(q76),
    .q77(q77),
    .q78(q78),
    .q81(q81),
    .q82(q82),
    .q83(q83),
    .q84(q84),
    .q85(q85),
    .q86(q86),
    .q87(q87),
    .q88(q88),
    .enable(valid_quan),
	.sram_waddr(sramB_waddr),
	.sram_wdata(sramB_wdata),
	.wen(sramB_wen),
	.valid(valid_RLC)
);

huffman U0(
    .clk(clk),
    .rst_n(rst_n),
    .valid(valid_RLC),
    .sram_data(sramB_rdata),
    .sram_addr(sramB_raddr),
    .code_length1(code_length1),
    .code_out1(code_out1),
    .code_length2(code_length2),
    .code_out2(code_out2),
    .code_length3(code_length3),
    .code_out3(code_out3),
    .code_length4(code_length4),
    .code_out4(code_out4),
    .code_length5(code_length5),
    .code_out5(code_out5),
    .code_length6(code_length6),
    .code_out6(code_out6),
    .code_length7(code_length7),
    .code_out7(code_out7),
    .code_length8(code_length8),
    .code_out8(code_out8),

    .code_length_DC(code_length_DC),
    .code_out_DC(code_out_DC),

    .code_length_table(code_length_table),
    .code_out_table(code_out_table),
    .out_valid(out_valid)
);


endmodule
